library verilog;
use verilog.vl_types.all;
entity lab2_2 is
    port(
        i               : in     vl_logic;
        s1              : in     vl_logic;
        s0              : in     vl_logic;
        y3              : out    vl_logic;
        y2              : out    vl_logic;
        y1              : out    vl_logic;
        y0              : out    vl_logic
    );
end lab2_2;
