library verilog;
use verilog.vl_types.all;
entity lab2_1 is
    port(
        Y0              : out    vl_logic;
        S1              : in     vl_logic;
        S0              : in     vl_logic;
        I               : in     vl_logic;
        Y1              : out    vl_logic;
        Y2              : out    vl_logic;
        Y3              : out    vl_logic
    );
end lab2_1;
