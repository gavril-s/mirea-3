library verilog;
use verilog.vl_types.all;
entity lab2_2_vlg_sample_tst is
    port(
        i               : in     vl_logic;
        s0              : in     vl_logic;
        s1              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end lab2_2_vlg_sample_tst;
